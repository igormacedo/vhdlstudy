LIBRARY ieee;
USE ieee.STD_LOGIC_1164.all;
USE ieee.STD_LOGIC_ARITH.all;
--USE ieee.STD_LOGIC_SIGNED.all;
USE ieee.STD_LOGIC_UNSIGNED.all;

ENTITY ula IS
GENERIC(N : INTEGER := 4);

PORT(
	E : IN INTEGER RANGE 0 TO N-1;
	A : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
	B : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);

	S : OUT STD_LOGIC_VECTOR(2*N-1 DOWNTO 0)
);

END ENTITY;

ARCHITECTURE estrutura OF ula IS

SIGNAL aux : STD_LOGIC_VECTOR(N-1 DOWNTO 0);

BEGIN
	aux <= (OTHERS => '0');
	WITH E SELECT
		S <= 	aux & (A+B) WHEN 0,
					A*B WHEN 1,
					aux & (A XOR B) WHEN 2,
					aux & (A AND B) WHEN 3;
END ARCHITECTURE;
